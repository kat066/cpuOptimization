`include "mips_core.svh"

interface instruction_Queue_ifc ();
	logic [1 : 0] Valid_Ready[31 : 0];
	decoder_output_ifc instruction[31 : 0]();
	logic [31 : 0] source [31 : 0][1 : 0];
	logic [31 : 0] destination [31 : 0];
	logic [31 : 0] active_List_Index[31 : 0];


endinterface


module instruction_Queue (
	decoder_output_ifc.in decoded
	decoder_output_ifc.out out
)
instruction_Queue_ifc Instr_Queue();
always_comb begin
	int count = 0;
	while (count < 32) begin

end


endmodule
