`include "mips_core.svh"
/* priority_encoder.sv
 *
 * Author: Haaris Tahir-Kheli
 * Date  : June 2nd, 2021
 *
 * A priority encoder that takes, as parameters, the number of inputs, 
 * and a wire signal to determine whether or not the encoder will operate
 * as a high priority encoder, or a low priority encoder.
 *
 * The output of the encoder is the binary encoding of the "index" of the
 * valid input that has the highest priority (based on whatever priority scheme the
 * module is uses, which is based on the value of the parameter, "HIGH_PRIORITY", 
 * and whether or not a 1 or a 0 is going to be seen as the valid input, which is
 * based on the value of the parameter, "SIGNAL".)
 * 
 */
module priority_encoder_64 #(parameter HIGH_PRIORITY = 0, parameter SIGNAL = 1) (
	input data_inputs[63:0],
	output logic [5:0] encoding_output
);

int i;

always_comb begin
	encoding_output = 0;
	
	if (HIGH_PRIORITY) begin
		for (int i = 0; i < 64; i++) begin
			if(data_inputs[i] == SIGNAL) begin
				encoding_output = i;
				break;
			end
		end	
	end
	else begin
		for (int i = 63; i >= 0; i--) begin
			if(data_inputs[i] == SIGNAL) begin
				encoding_output = i;
				break;
			end
		end		
	end


	/*
	packed_data_inputs[63:0] = { << {data_inputs[63:0]}};
	if (HIGH_PRIORITY) begin
		if (SIGNAL) begin
			casex(packed_data_inputs)
				64'b1XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd63;
				64'b01XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd62;
				64'b001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd61;
				64'b0001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd60;
				64'b00001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd59;
				64'b000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd58;
				64'b0000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd57;
				64'b00000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd56;
				64'b000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd55;
				64'b0000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd54;
				64'b00000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd53;
				64'b000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd52;
				64'b0000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd51;
				64'b00000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd50;
				64'b000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd49;
				64'b0000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd48;
				64'b00000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd47;
				64'b000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd46;
				64'b0000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd45;
				64'b00000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd44;
				64'b000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd43;
				64'b0000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd42;
				64'b00000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd41;
				64'b000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd40;
				64'b0000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd39;
				64'b00000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd38;
				64'b000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd37;
				64'b0000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd36;
				64'b00000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd35;
				64'b000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd34;
				64'b0000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd33;
				64'b00000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd32;
				64'b000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd31;
				64'b0000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd30;
				64'b00000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd29;
				64'b000000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd28;
				64'b0000000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd27;
				64'b00000000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd26;
				64'b000000000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd25;
				64'b0000000000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd24;
				64'b00000000000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd23;
				64'b000000000000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd22;
				64'b0000000000000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd21;
				64'b00000000000000000000000000000000000000000001XXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd20;	
				64'b000000000000000000000000000000000000000000001XXXXXXXXXXXXXXXXXXX: encoding_output = 6'd19;
				64'b0000000000000000000000000000000000000000000001XXXXXXXXXXXXXXXXXX: encoding_output = 6'd18;
				64'b00000000000000000000000000000000000000000000001XXXXXXXXXXXXXXXXX: encoding_output = 6'd17;
				64'b000000000000000000000000000000000000000000000001XXXXXXXXXXXXXXXX: encoding_output = 6'd16;
				64'b0000000000000000000000000000000000000000000000001XXXXXXXXXXXXXXX: encoding_output = 6'd15;
				64'b00000000000000000000000000000000000000000000000001XXXXXXXXXXXXXX: encoding_output = 6'd14;
				64'b000000000000000000000000000000000000000000000000001XXXXXXXXXXXXX: encoding_output = 6'd13;
				64'b0000000000000000000000000000000000000000000000000001XXXXXXXXXXXX: encoding_output = 6'd12;
				64'b00000000000000000000000000000000000000000000000000001XXXXXXXXXXX: encoding_output = 6'd11;
				64'b000000000000000000000000000000000000000000000000000001XXXXXXXXXX: encoding_output = 6'd10;
				64'b0000000000000000000000000000000000000000000000000000001XXXXXXXXX: encoding_output = 6'd9;
				64'b00000000000000000000000000000000000000000000000000000001XXXXXXXX: encoding_output = 6'd8;
				64'b000000000000000000000000000000000000000000000000000000001XXXXXXX: encoding_output = 6'd7;
				64'b0000000000000000000000000000000000000000000000000000000001XXXXXX: encoding_output = 6'd6;
				64'b00000000000000000000000000000000000000000000000000000000001XXXXX: encoding_output = 6'd5;
				64'b000000000000000000000000000000000000000000000000000000000001XXXX: encoding_output = 6'd4;
				64'b0000000000000000000000000000000000000000000000000000000000001XXX: encoding_output = 6'd3;
				64'b00000000000000000000000000000000000000000000000000000000000001XX: encoding_output = 6'd2;
				64'b000000000000000000000000000000000000000000000000000000000000001X: encoding_output = 6'd1;
				64'b0000000000000000000000000000000000000000000000000000000000000001: encoding_output = 6'd0;
				default																: encoding_output = 6'd0;
			endcase
		end
		else begin
			casex(packed_data_inputs)
				64'b0XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd63;
				64'b10XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd62;
				64'b110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd61;
				64'b1110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd60;
				64'b11110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd59;
				64'b111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd58;
				64'b1111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd57;
				64'b11111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd56;
				64'b111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd55;
				64'b1111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd54;
				64'b11111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd53;
				64'b111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd52;
				64'b1111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd51;
				64'b11111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd50;
				64'b111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd49;
				64'b1111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd48;
				64'b11111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd47;
				64'b111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd46;
				64'b1111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd45;
				64'b11111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd44;
				64'b111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd43;
				64'b1111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd42;
				64'b11111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd41;
				64'b111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd40;
				64'b1111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd39;
				64'b11111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd38;
				64'b111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd37;
				64'b1111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd36;
				64'b11111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd35;
				64'b111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd34;
				64'b1111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd33;
				64'b11111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd32;
				64'b111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd31;
				64'b1111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd30;
				64'b11111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd29;
				64'b111111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd28;
				64'b1111111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd27;
				64'b11111111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd26;
				64'b111111111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd25;
				64'b1111111111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd24;
				64'b11111111111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd23;
				64'b111111111111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd22;
				64'b1111111111111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd21;
				64'b11111111111111111111111111111111111111111110XXXXXXXXXXXXXXXXXXXX: encoding_output = 6'd20;	
				64'b111111111111111111111111111111111111111111110XXXXXXXXXXXXXXXXXXX: encoding_output = 6'd19;
				64'b1111111111111111111111111111111111111111111110XXXXXXXXXXXXXXXXXX: encoding_output = 6'd18;
				64'b11111111111111111111111111111111111111111111110XXXXXXXXXXXXXXXXX: encoding_output = 6'd17;
				64'b111111111111111111111111111111111111111111111110XXXXXXXXXXXXXXXX: encoding_output = 6'd16;
				64'b1111111111111111111111111111111111111111111111110XXXXXXXXXXXXXXX: encoding_output = 6'd15;
				64'b11111111111111111111111111111111111111111111111110XXXXXXXXXXXXXX: encoding_output = 6'd14;
				64'b111111111111111111111111111111111111111111111111110XXXXXXXXXXXXX: encoding_output = 6'd13;
				64'b1111111111111111111111111111111111111111111111111110XXXXXXXXXXXX: encoding_output = 6'd12;
				64'b11111111111111111111111111111111111111111111111111110XXXXXXXXXXX: encoding_output = 6'd11;
				64'b111111111111111111111111111111111111111111111111111110XXXXXXXXXX: encoding_output = 6'd10;
				64'b1111111111111111111111111111111111111111111111111111110XXXXXXXXX: encoding_output = 6'd9;
				64'b11111111111111111111111111111111111111111111111111111110XXXXXXXX: encoding_output = 6'd8;
				64'b111111111111111111111111111111111111111111111111111111110XXXXXXX: encoding_output = 6'd7;
				64'b1111111111111111111111111111111111111111111111111111111110XXXXXX: encoding_output = 6'd6;
				64'b11111111111111111111111111111111111111111111111111111111110XXXXX: encoding_output = 6'd5;
				64'b111111111111111111111111111111111111111111111111111111111110XXXX: encoding_output = 6'd4;
				64'b1111111111111111111111111111111111111111111111111111111111110XXX: encoding_output = 6'd3;
				64'b11111111111111111111111111111111111111111111111111111111111110XX: encoding_output = 6'd2;
				64'b111111111111111111111111111111111111111111111111111111111111110X: encoding_output = 6'd1;
				64'b1111111111111111111111111111111111111111111111111111111111111110: encoding_output = 6'd0;	
				default																: encoding_output = 6'd0;				
			endcase
		end
	end
	else begin
		if (SIGNAL) begin
			casex(packed_data_inputs)
				64'b1000000000000000000000000000000000000000000000000000000000000000: encoding_output = 6'd63;
				64'bX100000000000000000000000000000000000000000000000000000000000000: encoding_output = 6'd62;
				64'bXX10000000000000000000000000000000000000000000000000000000000000: encoding_output = 6'd61;
				64'bXXX1000000000000000000000000000000000000000000000000000000000000: encoding_output = 6'd60;
				64'bXXXX100000000000000000000000000000000000000000000000000000000000: encoding_output = 6'd59;
				64'bXXXXX10000000000000000000000000000000000000000000000000000000000: encoding_output = 6'd58;
				64'bXXXXXX1000000000000000000000000000000000000000000000000000000000: encoding_output = 6'd57;
				64'bXXXXXXX100000000000000000000000000000000000000000000000000000000: encoding_output = 6'd56;
				64'bXXXXXXXX10000000000000000000000000000000000000000000000000000000: encoding_output = 6'd55;
				64'bXXXXXXXXX1000000000000000000000000000000000000000000000000000000: encoding_output = 6'd54;
				64'bXXXXXXXXXX100000000000000000000000000000000000000000000000000000: encoding_output = 6'd53;
				64'bXXXXXXXXXXX10000000000000000000000000000000000000000000000000000: encoding_output = 6'd52;
				64'bXXXXXXXXXXXX1000000000000000000000000000000000000000000000000000: encoding_output = 6'd51;
				64'bXXXXXXXXXXXXX100000000000000000000000000000000000000000000000000: encoding_output = 6'd50;
				64'bXXXXXXXXXXXXXX10000000000000000000000000000000000000000000000000: encoding_output = 6'd49;
				64'bXXXXXXXXXXXXXXX1000000000000000000000000000000000000000000000000: encoding_output = 6'd48;
				64'bXXXXXXXXXXXXXXXX100000000000000000000000000000000000000000000000: encoding_output = 6'd47;
				64'bXXXXXXXXXXXXXXXXX10000000000000000000000000000000000000000000000: encoding_output = 6'd46;
				64'bXXXXXXXXXXXXXXXXXX1000000000000000000000000000000000000000000000: encoding_output = 6'd45;
				64'bXXXXXXXXXXXXXXXXXXX100000000000000000000000000000000000000000000: encoding_output = 6'd44;
				64'bXXXXXXXXXXXXXXXXXXXX10000000000000000000000000000000000000000000: encoding_output = 6'd43;
				64'bXXXXXXXXXXXXXXXXXXXXX1000000000000000000000000000000000000000000: encoding_output = 6'd42;
				64'bXXXXXXXXXXXXXXXXXXXXXX100000000000000000000000000000000000000000: encoding_output = 6'd41;
				64'bXXXXXXXXXXXXXXXXXXXXXXX10000000000000000000000000000000000000000: encoding_output = 6'd40;
				64'bXXXXXXXXXXXXXXXXXXXXXXXX1000000000000000000000000000000000000000: encoding_output = 6'd39;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXX100000000000000000000000000000000000000: encoding_output = 6'd38;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXX10000000000000000000000000000000000000: encoding_output = 6'd37;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXX1000000000000000000000000000000000000: encoding_output = 6'd36;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX100000000000000000000000000000000000: encoding_output = 6'd35;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10000000000000000000000000000000000: encoding_output = 6'd34;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000000000000000000000000000000000: encoding_output = 6'd33;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX100000000000000000000000000000000: encoding_output = 6'd32;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10000000000000000000000000000000: encoding_output = 6'd31;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000000000000000000000000000000: encoding_output = 6'd30;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX100000000000000000000000000000: encoding_output = 6'd29;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10000000000000000000000000000: encoding_output = 6'd28;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000000000000000000000000000: encoding_output = 6'd27;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX100000000000000000000000000: encoding_output = 6'd26;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10000000000000000000000000: encoding_output = 6'd25;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000000000000000000000000: encoding_output = 6'd24;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX100000000000000000000000: encoding_output = 6'd23;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10000000000000000000000: encoding_output = 6'd22;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000000000000000000000: encoding_output = 6'd21;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX100000000000000000000: encoding_output = 6'd20;	
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10000000000000000000: encoding_output = 6'd19;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000000000000000000: encoding_output = 6'd18;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX100000000000000000: encoding_output = 6'd17;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10000000000000000: encoding_output = 6'd16;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000000000000000: encoding_output = 6'd15;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX100000000000000: encoding_output = 6'd14;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10000000000000: encoding_output = 6'd13;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000000000000: encoding_output = 6'd12;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX100000000000: encoding_output = 6'd11;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10000000000: encoding_output = 6'd10;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000000000: encoding_output = 6'd9;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX100000000: encoding_output = 6'd8;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10000000: encoding_output = 6'd7;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000000: encoding_output = 6'd6;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX100000: encoding_output = 6'd5;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10000: encoding_output = 6'd4;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000: encoding_output = 6'd3;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX100: encoding_output = 6'd2;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10: encoding_output = 6'd1;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1: encoding_output = 6'd0;	
				default																: encoding_output = 6'd0;				
			endcase	
		end
		else begin
			casex(packed_data_inputs)
				64'b0111111111111111111111111111111111111111111111111111111111111111: encoding_output = 6'd63;
				64'bX011111111111111111111111111111111111111111111111111111111111111: encoding_output = 6'd62;
				64'bXX01111111111111111111111111111111111111111111111111111111111111: encoding_output = 6'd61;
				64'bXXX0111111111111111111111111111111111111111111111111111111111111: encoding_output = 6'd60;
				64'bXXXX011111111111111111111111111111111111111111111111111111111111: encoding_output = 6'd59;
				64'bXXXXX01111111111111111111111111111111111111111111111111111111111: encoding_output = 6'd58;
				64'bXXXXXX0111111111111111111111111111111111111111111111111111111111: encoding_output = 6'd57;
				64'bXXXXXXX011111111111111111111111111111111111111111111111111111111: encoding_output = 6'd56;
				64'bXXXXXXXX01111111111111111111111111111111111111111111111111111111: encoding_output = 6'd55;
				64'bXXXXXXXXX0111111111111111111111111111111111111111111111111111111: encoding_output = 6'd54;
				64'bXXXXXXXXXX011111111111111111111111111111111111111111111111111111: encoding_output = 6'd53;
				64'bXXXXXXXXXXX01111111111111111111111111111111111111111111111111111: encoding_output = 6'd52;
				64'bXXXXXXXXXXXX0111111111111111111111111111111111111111111111111111: encoding_output = 6'd51;
				64'bXXXXXXXXXXXXX011111111111111111111111111111111111111111111111111: encoding_output = 6'd50;
				64'bXXXXXXXXXXXXXX01111111111111111111111111111111111111111111111111: encoding_output = 6'd49;
				64'bXXXXXXXXXXXXXXX0111111111111111111111111111111111111111111111111: encoding_output = 6'd48;
				64'bXXXXXXXXXXXXXXXX011111111111111111111111111111111111111111111111: encoding_output = 6'd47;
				64'bXXXXXXXXXXXXXXXXX01111111111111111111111111111111111111111111111: encoding_output = 6'd46;
				64'bXXXXXXXXXXXXXXXXXX0111111111111111111111111111111111111111111111: encoding_output = 6'd45;
				64'bXXXXXXXXXXXXXXXXXXX011111111111111111111111111111111111111111111: encoding_output = 6'd44;
				64'bXXXXXXXXXXXXXXXXXXXX01111111111111111111111111111111111111111111: encoding_output = 6'd43;
				64'bXXXXXXXXXXXXXXXXXXXXX0111111111111111111111111111111111111111111: encoding_output = 6'd42;
				64'bXXXXXXXXXXXXXXXXXXXXXX011111111111111111111111111111111111111111: encoding_output = 6'd41;
				64'bXXXXXXXXXXXXXXXXXXXXXXX01111111111111111111111111111111111111111: encoding_output = 6'd40;
				64'bXXXXXXXXXXXXXXXXXXXXXXXX0111111111111111111111111111111111111111: encoding_output = 6'd39;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXX011111111111111111111111111111111111111: encoding_output = 6'd38;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXX01111111111111111111111111111111111111: encoding_output = 6'd37;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXX0111111111111111111111111111111111111: encoding_output = 6'd36;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX011111111111111111111111111111111111: encoding_output = 6'd35;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01111111111111111111111111111111111: encoding_output = 6'd34;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111111111111111111111111111111111: encoding_output = 6'd33;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX011111111111111111111111111111111: encoding_output = 6'd32;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01111111111111111111111111111111: encoding_output = 6'd31;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111111111111111111111111111111: encoding_output = 6'd30;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX011111111111111111111111111111: encoding_output = 6'd29;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01111111111111111111111111111: encoding_output = 6'd28;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111111111111111111111111111: encoding_output = 6'd27;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX011111111111111111111111111: encoding_output = 6'd26;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01111111111111111111111111: encoding_output = 6'd25;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111111111111111111111111: encoding_output = 6'd24;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX011111111111111111111111: encoding_output = 6'd23;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01111111111111111111111: encoding_output = 6'd22;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111111111111111111111: encoding_output = 6'd21;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX011111111111111111111: encoding_output = 6'd20;	
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01111111111111111111: encoding_output = 6'd19;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111111111111111111: encoding_output = 6'd18;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX011111111111111111: encoding_output = 6'd17;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01111111111111111: encoding_output = 6'd16;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111111111111111: encoding_output = 6'd15;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX011111111111111: encoding_output = 6'd14;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01111111111111: encoding_output = 6'd13;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111111111111: encoding_output = 6'd12;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX011111111111: encoding_output = 6'd11;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01111111111: encoding_output = 6'd10;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111111111: encoding_output = 6'd9;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX011111111: encoding_output = 6'd8;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01111111: encoding_output = 6'd7;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111111: encoding_output = 6'd6;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX011111: encoding_output = 6'd5;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01111: encoding_output = 6'd4;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111: encoding_output = 6'd3;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX011: encoding_output = 6'd2;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX01: encoding_output = 6'd1;
				64'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0: encoding_output = 6'd0;	
				default																: encoding_output = 6'd0;				
			endcase			
		end
	end
	*/
end

endmodule
