`include "mips_core.svh"


module free_List(
	
);

logic free [64];
always_comb begin
	int count = 0;
	while (count < 32) begin

	end

end
endmodule

